package nn_param_pkg;

  localparam INT_BITS  = 6;
  localparam FRC_BITS  = 7;
  localparam BITS      = 13;
  
  localparam PICT_SIZE = 28;
  localparam WIDTH     = 784;

  localparam ADDR_RC   = 5;
  localparam ADDR_OUT  = 10;

  localparam RCO_TYPE  = 2;

  localparam NN_FSM_BUS_WIDTH  = 5;
    
endpackage